set_property -dict { PACKAGE_PIN U7   IOSTANDARD LVCMOS33 } [get_ports {num[0]}]
set_property -dict { PACKAGE_PIN V5   IOSTANDARD LVCMOS33 } [get_ports {num[1]}]
set_property -dict { PACKAGE_PIN U5   IOSTANDARD LVCMOS33 } [get_ports {num[2]}]
set_property -dict { PACKAGE_PIN V8   IOSTANDARD LVCMOS33 } [get_ports {num[3]}]
set_property -dict { PACKAGE_PIN U8   IOSTANDARD LVCMOS33 } [get_ports {num[4]}]
set_property -dict { PACKAGE_PIN W6   IOSTANDARD LVCMOS33 } [get_ports {num[5]}]
set_property -dict { PACKAGE_PIN W7   IOSTANDARD LVCMOS33 } [get_ports {num[6]}]
set_property -dict { PACKAGE_PIN V7   IOSTANDARD LVCMOS33 } [get_ports {num[7]}]

set_property PACKAGE_PIN W5 [get_ports Clk]							
	set_property IOSTANDARD LVCMOS33 [get_ports Clk]
	create_clock -add -name sys_clk_pin -period 10.00 -waveform {0 5} [get_ports Clk]

set_property PACKAGE_PIN V17 [get_ports {EIN}]					
	set_property IOSTANDARD LVCMOS33 [get_ports {EIN}]
set_property PACKAGE_PIN T17 [get_ports {RST}]					
	set_property IOSTANDARD LVCMOS33 [get_ports {RST}]
set_property PACKAGE_PIN W19 [get_ports {Submit}]					
	set_property IOSTANDARD LVCMOS33 [get_ports {Submit}]
set_property PACKAGE_PIN R2 [get_ports {rigged_win}]					
	set_property IOSTANDARD LVCMOS33 [get_ports {rigged_win}]
set_property PACKAGE_PIN T1 [get_ports {rigged_lose}]					
	set_property IOSTANDARD LVCMOS33 [get_ports {rigged_lose}]

set_property PACKAGE_PIN U2 [get_ports {anodes[0]}]					
	set_property IOSTANDARD LVCMOS33 [get_ports {anodes[0]}]
set_property PACKAGE_PIN U4 [get_ports {anodes[1]}]					
	set_property IOSTANDARD LVCMOS33 [get_ports {anodes[1]}]
set_property PACKAGE_PIN V4 [get_ports {anodes[2]}]					
	set_property IOSTANDARD LVCMOS33 [get_ports {anodes[2]}]
set_property PACKAGE_PIN W4 [get_ports {anodes[3]}]					
	set_property IOSTANDARD LVCMOS33 [get_ports {anodes[3]}]
